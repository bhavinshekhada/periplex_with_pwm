`define TOTAL_UART 1
`define TOTAL_GPIO_CTRLS 1
`define TOTAL_PWM 3
`define TOTAL_I2C 0
    